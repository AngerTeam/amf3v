module amf3v

const amf_undefined := 0
const amf_null := 1
const amf_false := 2
const amf_true := 3
const amf_packed_int := 4
const amf_double := 5
const amf_string := 6
const amf_xml_object := 7
const amf_date := 8
const amf_array := 9
const amf_object := 10
const amf_xml := 11
const amf_byte_array := 12
