module amf3v

pub struct AmfObject {

}
